grammar edu:umn:cs:melt:exts:ableC:halide:src;

exports edu:umn:cs:melt:exts:ableC:halide:src:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:halide:src:concretesyntax;

