grammar edu:umn:cs:melt:exts:ableC:halide;

exports edu:umn:cs:melt:exts:ableC:halide:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:halide:concretesyntax;

