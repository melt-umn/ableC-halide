grammar edu:umn:cs:melt:exts:ableC:halide:abstractsyntax;

imports silver:langutil;
imports silver:langutil:pp;
imports core:monad;

imports edu:umn:cs:melt:ableC:abstractsyntax:host;
imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:overloadable;
imports edu:umn:cs:melt:ableC:abstractsyntax:env;

global builtin::Location = builtinLoc("halide");

abstract production transformStmt
top::Stmt ::= s::Stmt t::Transformation
{
  top.pp =
    ppConcat([pp"transform ", braces(nestlines(2, s.pp)), pp" by ", braces(nestlines(2, t.pp))]);
  top.functionDefs := [];
  
  local normalizedS::Stmt = s.normalizeLoops.fromJust;
  normalizedS.env = s.env;
  normalizedS.returnType = s.returnType;
  
  t.iterStmtIn = stmtToIterStmt(normalizedS);
  
  local transResult::IterStmt = t.iterStmtOut;
  transResult.env = top.env;
  transResult.returnType = top.returnType;
  
  forwards to unsafeTrace(
    if !null(s.errors)
    then warnStmt(s.errors)
    else if !null(t.errors)
    then warnStmt(t.errors)
    else if !null(normalizedS.errors)
    then warnStmt(normalizedS.errors) -- Shouldn't happen
    else if !null(transResult.errors)
    then warnStmt(transResult.errors) -- Shouldn't happen
    else transResult.hostTrans,
    print(hackUnparse(normalizedS), unsafeIO()));
}

function isSimple
Boolean ::= e::Expr
{
  -- Avoid decorating with the full env during rewriting.
  -- This will never make an otherwise-not-simple AST appear simple.
  e.env = emptyEnv();
  e.returnType = nothing();
  return e.isSimple;
}

function isIntConst
Boolean ::= e::Expr
{
  -- Avoid decorating with the full env during rewriting.
  -- This will never make an non-int-constant AST appear to be an int constant.
  e.env = emptyEnv();
  e.returnType = nothing();
  return e.integerConstantValue.isJust;
}

function intValue
Integer ::= e::Expr
{
  -- Avoid decorating with the full env during rewriting.
  -- This will never make an non-int-constant AST appear to be an int constant.
  e.env = emptyEnv();
  e.returnType = nothing();
  return e.integerConstantValue.fromJust;
}

strategy attribute simplifyNumericExprStep =
  rule on Expr of
  -- Simplify expressions as much as possible
  | ableC_Expr { ($Expr{e}) } -> e
  | ableC_Expr { -$Expr{e} } when isIntConst(e) -> mkIntConst(-intValue(e), builtin)
  | ableC_Expr { $Expr{e1} + $Expr{e2} } when isIntConst(e1) && isIntConst(e2) ->
    mkIntConst(intValue(e1) + intValue(e2), builtin)
  | ableC_Expr { $Expr{e1} - $Expr{e2} } when isIntConst(e1) && isIntConst(e2) ->
    mkIntConst(intValue(e1) - intValue(e2), builtin)
  | ableC_Expr { $Expr{e1} * $Expr{e2} } when isIntConst(e1) && isIntConst(e2) ->
    mkIntConst(intValue(e1) * intValue(e2), builtin)
  | ableC_Expr { $Expr{e1} / $Expr{e2} } when isIntConst(e1) && isIntConst(e2) && intValue(e2) > 0 ->
    mkIntConst(intValue(e1) / intValue(e2), builtin)
  end;

strategy attribute simplifyNumericExpr = innermost(simplifyNumericExprStep);
strategy attribute simplifyLoopExprs =
  forDeclStmt(simplifyNumericExpr, simplifyNumericExpr, simplifyNumericExpr, id);

attribute simplifyNumericExprStep, simplifyNumericExpr, simplifyLoopExprs occurs on
  Stmt, Decl, Declarators, Declarator, MaybeInitializer, Initializer, MaybeExpr, Expr;
propagate simplifyNumericExprStep, simplifyNumericExpr, simplifyLoopExprs on
  Stmt, Decl, Declarators, Declarator, MaybeInitializer, Initializer, MaybeExpr, Expr;

strategy attribute preprocessLoop =
  rule on Stmt of
  -- Normalize condition orderings
  | ableC_Stmt { for ($BaseTypeExpr{t} $Name{i1} = $Expr{initial}; $Expr{limit} < $Name{i2}; $Expr{iter}) $Stmt{b} }
      when i1.name == i2.name ->
    ableC_Stmt { for ($BaseTypeExpr{t} $Name{i1} = $Expr{initial}; $Name{i2} > $Expr{limit}; $Expr{iter}) $Stmt{b} }
  | ableC_Stmt { for ($BaseTypeExpr{t} $Name{i1} = $Expr{initial}; $Expr{limit} > $Name{i2}; $Expr{iter}) $Stmt{b} }
      when i1.name == i2.name ->
    ableC_Stmt { for ($BaseTypeExpr{t} $Name{i1} = $Expr{initial}; $Name{i2} < $Expr{limit}; $Expr{iter}) $Stmt{b} }
  | ableC_Stmt { for ($BaseTypeExpr{t} $Name{i1} = $Expr{initial}; $Expr{limit} <= $Name{i2}; $Expr{iter}) $Stmt{b} }
      when i1.name == i2.name ->
    ableC_Stmt { for ($BaseTypeExpr{t} $Name{i1} = $Expr{initial}; $Name{i2} >= $Expr{limit}; $Expr{iter}) $Stmt{b} }
  | ableC_Stmt { for ($BaseTypeExpr{t} $Name{i1} = $Expr{initial}; $Expr{limit} >= $Name{i2}; $Expr{iter}) $Stmt{b} }
      when i1.name == i2.name ->
    ableC_Stmt { for ($BaseTypeExpr{t} $Name{i1} = $Expr{initial}; $Name{i2} <= $Expr{limit}; $Expr{iter}) $Stmt{b} }
  
  -- Normalize condition operators
  | ableC_Stmt { for ($Decl{init} $Name{i} <= $Expr{limit}; $Expr{iter}) $Stmt{b} } ->
    ableC_Stmt { for ($Decl{init} $Name{i} < $Expr{limit} + 1; $Expr{iter}) $Stmt{b} }
  | ableC_Stmt { for ($Decl{init} $Name{i} > $Expr{limit}; $Expr{iter}) $Stmt{b} } ->
    ableC_Stmt { for ($Decl{init} $Name{i} >= $Expr{limit} + 1; $Expr{iter}) $Stmt{b} }
  
  -- Expand increment/decrement operators
  | ableC_Stmt { for ($Decl{init} $Expr{cond}; $Name{i}++) $Stmt{b} } ->
    ableC_Stmt { for ($Decl{init} $Expr{cond}; $Name{i} += 1) $Stmt{b} }
  | ableC_Stmt { for ($Decl{init} $Expr{cond}; $Name{i}--) $Stmt{b} } ->
    ableC_Stmt { for ($Decl{init} $Expr{cond}; $Name{i} -= 1) $Stmt{b} }
  end;

-- Functor transformation to perform a renaming over anything
-- Not capture-avoiding, but that's OK!
-- If we rename a shadowed name, then we will also rename the shadowing declaration.
autocopy attribute targetName::String;
autocopy attribute replacement::String;
functor attribute renamed;
aspect production name
top::Name ::= n::String
{
  top.renamed =
    if n == top.targetName
    then name(top.replacement, location=top.location)
    else top;
}

attribute targetName, replacement, renamed occurs on
  Name, MaybeName,
  GlobalDecls, Decls, Decl, Declarators, Declarator, FunctionDecl, Parameters, ParameterDecl, StructDecl, UnionDecl, EnumDecl, StructItemList, EnumItemList, StructItem, StructDeclarators, StructDeclarator, EnumItem,
  MemberDesignator,
  Expr, GenericAssocs, GenericAssoc,
  TypeName, BaseTypeExpr, TypeModifierExpr, TypeNames,
  NumericConstant,
  MaybeExpr, Exprs, ExprOrTypeName,
  Stmt,
  MaybeInitializer, Initializer, InitList, Init, Designator,
  SpecialSpecifiers;
propagate renamed on
  Name, MaybeName,
  GlobalDecls, Decls, Decl, Declarators, Declarator, FunctionDecl, Parameters, ParameterDecl, StructDecl, UnionDecl, EnumDecl, StructItemList, EnumItemList, StructItem, StructDeclarators, StructDeclarator, EnumItem,
  MemberDesignator,
  Expr, GenericAssocs, GenericAssoc,
  TypeName, BaseTypeExpr, TypeModifierExpr, TypeNames,
  NumericConstant,
  MaybeExpr, Exprs, ExprOrTypeName,
  Stmt,
  MaybeInitializer, Initializer, InitList, Init, Designator,
  SpecialSpecifiers
  excluding name;

aspect production forDeclStmt
top::Stmt ::= i::Decl  c::MaybeExpr  s::MaybeExpr  b::Stmt
{
  local iName::String =
    case i of
    | ableC_Decl { $BaseTypeExpr{_} $Name{name(n)} = $Expr{_}; } -> n
    | _ -> error("Only should be demanded for a variable initializer")
    end;
  b.targetName = iName;
  b.replacement = s"_iter_${iName}_${toString(genInt())}";
}

strategy attribute transLoop =
  rule on Stmt of
  -- Restore increment operator on loops that are otherwise-normal
  | ableC_Stmt {
      for ($BaseTypeExpr{t} $Name{i1} = 0; $Name{i2} < $Expr{n}; $Name{i3} += 1) $Stmt{b}
    } when i1.name == i2.name && i1.name == i3.name ->
    ableC_Stmt {
      for ($BaseTypeExpr{t} $Name{i1} = 0; $Name{i2} < $Expr{n}; $Name{i3}++) $Stmt{b}
    }
  
  -- Normalize loops with nonstandard initial or step values
  | ableC_Stmt {
      for ($BaseTypeExpr{t} $Name{i1} = $Expr{initial}; $Name{i2} < $Expr{limit}; $Name{i3} += $Expr{step})
        $Stmt{b}
    } when i1.name == i2.name && i1.name == i3.name && isSimple(initial) && isSimple(step) ->
      ableC_Stmt {
        for ($BaseTypeExpr{t} $Name{i1} = 0; $Name{i2} < ($Expr{limit} - $Expr{initial}) / $Expr{step}; $Name{i3}++) {
          typeof($Name{i1}) $name{b.replacement} = $Expr{initial} + $Name{i1} * $Expr{step};
          $Stmt{b.renamed}
        }
      }
  
  -- Normalize "backwards" loops, possibly with with nonstandard initial or step values
  | ableC_Stmt {
      for ($BaseTypeExpr{t} $Name{i1} = $Expr{initial}; $Name{i2} >= $Expr{limit}; $Name{i3} -= $Expr{step})
        $Stmt{b}
    } when i1.name == i2.name && i1.name == i3.name && isSimple(initial) && isSimple(step) ->
      ableC_Stmt {
        for ($BaseTypeExpr{t} $Name{i1} = 0; $Name{i2} < ($Expr{initial} - $Expr{limit} + 1) / $Expr{step}; $Name{i3}++) {
          typeof($Name{i1}) $name{b.replacement} = $Expr{initial} - $Name{i1} * $Expr{step};
          $Stmt{b.renamed}
        }
      }
  end;

strategy attribute normalizeLoops =
  bottomUp(try(simplifyLoopExprs <* repeat(preprocessLoop))) <*
  topDown(try(transLoop <* simplifyLoopExprs));

attribute preprocessLoop, transLoop, normalizeLoops occurs on Stmt;
propagate preprocessLoop, transLoop, normalizeLoops on Stmt;

function stmtToIterStmt
IterStmt ::= s::Decorated Stmt
{
  return
    case s of
    | nullStmt() -> nullIterStmt()
    | seqStmt(s1, s2) -> seqIterStmt(stmtToIterStmt(s1), stmtToIterStmt(s2))
    | compoundStmt(s1) -> stmtToIterStmt(s1)
    | ableC_Stmt { if ($Expr{c}) $Stmt{t} else $Stmt{e} } ->
      condIterStmt(c, stmtToIterStmt(t), stmtToIterStmt(e))
    | ableC_Stmt {
        for ($BaseTypeExpr{t} $Name{i1} = 0; $Name{i2} host::< $Expr{n}; $Name{i3} host::++)
          $Stmt{b}
      } when i1.name == i2.name && i1.name == i3.name ->
      forIterStmt(t, baseTypeExpr(), i1, n, stmtToIterStmt(b))
    | s -> stmtIterStmt(new(s))
    end;
}

abstract production multiForStmt
top::Stmt ::= ivs::IterVars body::Stmt
{
  top.pp = pp"forall (${ivs.pp}) ${braces(nestlines(2, body.pp))}";
  top.functionDefs := [];
  
  ivs.forIterStmtBody = stmtIterStmt(body);
  forwards to ivs.forIterStmtTrans.hostTrans;
}

monoid attribute iterDefs::[Def] with [], ++;
synthesized attribute hostTrans::Stmt;

nonterminal IterStmt with pp, errors, defs, iterDefs, hostTrans, env, returnType;

propagate iterDefs on IterStmt;

abstract production nullIterStmt
top::IterStmt ::= 
{
  propagate errors, defs;
  top.pp = notext();
  top.hostTrans = nullStmt();
}

abstract production seqIterStmt
top::IterStmt ::= h::IterStmt t::IterStmt
{
  propagate errors, defs;
  top.pp = ppConcat([ h.pp, line(), t.pp ]);
  top.hostTrans = seqStmt(h.hostTrans, t.hostTrans);
  
  t.env = addEnv(h.defs, h.env);
}

abstract production compoundIterStmt
top::IterStmt ::= is::IterStmt
{
  propagate errors;
  top.pp = braces(nestlines(2, is.pp));
  top.defs := [];
  top.hostTrans = compoundStmt(is.hostTrans);
  
  is.env = openScopeEnv(top.env);
}

abstract production stmtIterStmt
top::IterStmt ::= s::Stmt
{
  propagate errors, defs;
  top.pp = braces(braces(nestlines(2, s.pp)));
  top.hostTrans = s;
}

abstract production condIterStmt
top::IterStmt ::= cond::Expr th::IterStmt el::IterStmt
{
  propagate errors, defs;
  top.pp = pp"if (${cond.pp})${nestlines(2, th.pp)} else ${nestlines(2, el.pp)}";
  top.hostTrans = ifStmt(cond, th.hostTrans, el.hostTrans);
}

abstract production forIterStmt
top::IterStmt ::= bty::BaseTypeExpr mty::TypeModifierExpr n::Name cutoff::Expr body::IterStmt
{
  top.pp = pp"for (${ppConcat([bty.pp, space(), mty.lpp, n.pp, mty.rpp])} : ${cutoff.pp}) ${braces(nestlines(2, body.pp))}";
  top.errors := bty.errors ++ d.errors ++ cutoff.errors ++ body.errors;
  top.errors <- n.valueRedeclarationCheckNoCompatible;
  
  production d::Declarator =
    declarator(
      n, mty, nilAttribute(),
      justInitializer(exprInitializer(ableC_Expr {0})));
  d.env = openScopeEnv(top.env);
  d.baseType = bty.typerep;
  d.typeModifierIn = bty.typeModifier;
  d.isTopLevel = false;
  d.isTypedef = false;
  d.givenStorageClasses = nilStorageClass();
  d.givenAttributes = nilAttribute();
  d.returnType = top.returnType;
  
  top.defs := [];
  top.iterDefs <- [valueDef(n.name, declaratorValueItem(d))];
  top.hostTrans =
    ableC_Stmt {
      for ($Decl{
        variableDecls(
          nilStorageClass(), nilAttribute(),
          bty,
          consDeclarator(d, nilDeclarator()))} $Name{n} < $Expr{cutoff}; $Name{n}++)
        $Stmt{body.hostTrans}
    };
  
  bty.givenRefId = nothing();
  body.env = addEnv(d.defs, openScopeEnv(top.env));
}

abstract production parallelForIterStmt
top::IterStmt ::= numThreads::Maybe<Integer> bty::BaseTypeExpr mty::TypeModifierExpr n::Name cutoff::Expr body::IterStmt
{
  local numThreadsPP::Document =
    case numThreads of
    | just(n) -> parens(text(toString(n)))
    | nothing() -> notext()
    end;
  top.pp = pp"for parallel${numThreadsPP} (${ppConcat([bty.pp, space(), mty.lpp, n.pp, mty.rpp])} : ${cutoff.pp}) ${braces(nestlines(2, body.pp))}";
  top.errors := bty.errors ++ d.errors ++ cutoff.errors ++ body.errors;
  top.errors <- n.valueRedeclarationCheckNoCompatible;
  
  production d::Declarator = declarator(n, mty, nilAttribute(), nothingInitializer());
  d.env = openScopeEnv(top.env);
  d.baseType = bty.typerep;
  d.typeModifierIn = bty.typeModifier;
  d.isTopLevel = false;
  d.isTypedef = false;
  d.givenStorageClasses = nilStorageClass();
  d.givenAttributes = nilAttribute();
  d.returnType = top.returnType;
  
  top.defs := [];
  
  {- TODO: We don't right now have a way to insert pragmas via abstract syntax, and OpenMP is
   - rather picky about the loop variable being declared in the loop and extra parentheses in the
   - predicate, so we need to resort to some hacks with txtStmt for now.
   -}
  top.hostTrans =
    compoundStmt(
      foldStmt([
        declStmt( -- Still re-declare the loop variable in the ast, so it shows up in env for the host error check
          variableDecls(
            nilStorageClass(), nilAttribute(),
            bty,
            consDeclarator(d, nilDeclarator()))),
        case numThreads of
          just(n) -> txtStmt(s"#pragma omp parallel for num_threads(${toString(n)})")
        | nothing() -> txtStmt("#pragma omp parallel for")
        end,
        txtStmt(s"for (${show(80, bty.pp)} ${show(80, head(d.pps))} = 0; ${n.name} < ${show(80, cutoff.pp)}; ${n.name}++)"),
        compoundStmt(body.hostTrans)]));
  
  bty.givenRefId = nothing();
  
  body.env = addEnv(d.defs, openScopeEnv(top.env));
}

abstract production vectorForIterStmt
top::IterStmt ::= bty::BaseTypeExpr mty::TypeModifierExpr n::Name cutoff::Expr body::IterStmt
{
  top.pp = pp"for vector (${ppConcat([bty.pp, space(), mty.lpp, n.pp, mty.rpp])} : ${cutoff.pp}) ${braces(nestlines(2, body.pp))}";
  top.errors := bty.errors ++ d.errors ++ cutoff.errors ++ body.errors;
  top.errors <- n.valueRedeclarationCheckNoCompatible;
  
  production d::Declarator = declarator(n, mty, nilAttribute(), nothingInitializer());
  d.env = openScopeEnv(top.env);
  d.baseType = bty.typerep;
  d.typeModifierIn = bty.typeModifier;
  d.isTopLevel = false;
  d.isTypedef = false;
  d.givenStorageClasses = nilStorageClass();
  d.givenAttributes = nilAttribute();
  d.returnType = top.returnType;
  
  top.defs := [];
  
  {- TODO: We don't right now have a way to insert pragmas via abstract syntax, and OpenMP is
   - rather picky about the loop variable being declared in the loop and extra parentheses in the
   - predicate, so we need to resort to some hacks with txtStmt for now.
   -}
  top.hostTrans =
    compoundStmt(
      foldStmt([
        declStmt( -- Still re-declare the loop variable in the ast, so it shows up in env for the host error check
          variableDecls(
            nilStorageClass(), nilAttribute(),
            bty,
            consDeclarator(d, nilDeclarator()))),
        txtStmt("#pragma omp simd"),
        txtStmt(s"for (${show(80, bty.pp)} ${show(80, head(d.pps))} = 0; ${n.name} < ${show(80, cutoff.pp)}; ${n.name}++)"),
        compoundStmt(body.hostTrans)]));
  
  bty.givenRefId = nothing();
  
  body.env = addEnv(d.defs, openScopeEnv(top.env));
}

synthesized attribute iterVarNames::[Name];

synthesized attribute forIterStmtTrans::IterStmt;
inherited attribute forIterStmtBody::IterStmt;

nonterminal IterVars with pp, errors, iterVarNames, forIterStmtTrans, forIterStmtBody, env, returnType;

propagate errors on IterVars;

abstract production consIterVar
top::IterVars ::= bty::BaseTypeExpr mty::TypeModifierExpr n::Name cutoff::Expr rest::IterVars
{
  top.pp = ppConcat([bty.pp, space(), mty.lpp, n.pp, mty.rpp, text(" : "), cutoff.pp, comma(), space(), rest.pp]);
  top.errors <-
    case cutoff.integerConstantValue of
    | just(n) when n < 1 -> [err(cutoff.location, "Split loop size must be >= 1")]
    | _ -> []
    end;
  top.iterVarNames = n :: rest.iterVarNames;
  
  top.forIterStmtTrans = forIterStmt(bty, mty, n, cutoff, rest.forIterStmtTrans);
  rest.forIterStmtBody = top.forIterStmtBody;
  
  bty.givenRefId = nothing();
  
  mty.baseType = bty.typerep;
  mty.typeModifierIn = bty.typeModifier;
}

abstract production consAnonIterVar
top::IterVars ::= cutoff::Expr rest::IterVars
{
  top.pp = ppConcat([cutoff.pp, comma(), rest.pp]);
  forwards to
    consIterVar(
      directTypeExpr(cutoff.typerep),
      baseTypeExpr(),
      name("_iter_var_" ++ toString(genInt()), location=builtin),
      cutoff, rest);
}

abstract production nilIterVar
top::IterVars ::= 
{
  top.pp = notext();
  top.iterVarNames = [];
  top.forIterStmtTrans = top.forIterStmtBody;
}

synthesized attribute iterVarName::Name;

inherited attribute forIterStmtCutoff::Expr;

nonterminal IterVar with pp, errors, iterVarName, forIterStmtTrans, forIterStmtCutoff, forIterStmtBody, env, returnType;

propagate errors on IterVar;

abstract production iterVar
top::IterVar ::= bty::BaseTypeExpr mty::TypeModifierExpr n::Name
{
  top.pp = ppConcat([bty.pp, space(), mty.lpp, n.pp, mty.rpp]);
  top.iterVarName = n;
  top.forIterStmtTrans = forIterStmt(bty, mty, n, top.forIterStmtCutoff, top.forIterStmtBody);
  
  bty.givenRefId = nothing();
  
  mty.baseType = bty.typerep;
  mty.typeModifierIn = bty.typeModifier;
}
